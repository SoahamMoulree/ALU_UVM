`define num_txns 200
`define W 8
`define N 4
`define SHIFT_WIDTH  $clog2(`W)

