class alu_seqr extends uvm_sequencer#(seq_item);

  `uvm_component_utils(alu_seqr)

  function new(string name,uvm_component parent);
    super.new(name,parent);
  endfunction

  endclass
