`include "uvm_macros.svh"
package alu_pkg;
  import uvm_pkg::*;
  `include "seq_item.sv"
  `include "sequence.sv"
  `include "sequencer.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "agent.sv"
  `include "scoreboard.sv"
  `include "coverage.sv"
  `include "environment.sv"
  `include "test.sv"
endpackage
